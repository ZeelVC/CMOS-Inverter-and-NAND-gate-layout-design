magic
tech scmos
timestamp 1734185267
<< nwell >>
rect -17 -10 17 36
<< ntransistor >>
rect -5 -42 -3 -32
rect 3 -42 5 -32
<< ptransistor >>
rect -5 -3 -3 17
rect 3 -3 5 17
<< ndiffusion >>
rect -6 -42 -5 -32
rect -3 -42 3 -32
rect 5 -41 6 -32
rect 5 -42 10 -41
<< pdiffusion >>
rect -6 -3 -5 17
rect -3 16 3 17
rect -3 -3 -2 16
rect 2 -3 3 16
rect 5 -2 6 17
rect 5 -3 10 -2
<< ndcontact >>
rect -10 -42 -6 -32
rect 6 -41 10 -32
<< pdcontact >>
rect -10 -3 -6 17
rect -2 -3 2 16
rect 6 -2 10 17
<< psubstratepcontact >>
rect -10 -50 -6 -46
rect -2 -50 2 -46
rect 6 -50 10 -46
<< nsubstratencontact >>
rect -10 28 -6 32
rect -2 28 2 32
rect 6 28 10 32
<< polysilicon >>
rect -5 17 -3 26
rect 3 17 5 26
rect -5 -32 -3 -3
rect 3 -32 5 -3
rect -5 -44 -3 -42
rect 3 -44 5 -42
<< polycontact >>
rect -9 -21 -5 -17
rect 5 -17 9 -13
<< metal1 >>
rect -6 28 -2 32
rect 2 28 6 32
rect -10 17 -6 28
rect 6 17 10 28
rect -14 -21 -9 -17
rect -2 -20 2 -3
rect 9 -17 15 -13
rect -2 -24 10 -20
rect 6 -32 10 -24
rect -10 -46 -6 -42
rect -6 -50 -2 -46
rect 2 -50 6 -46
<< labels >>
rlabel metal1 -4 30 -4 30 1 vdd
rlabel metal1 -4 -48 -4 -48 1 gnd
rlabel metal1 -12 -19 -12 -19 3 A
rlabel metal1 13 -15 13 -15 7 B
rlabel metal1 8 -22 8 -22 1 Y
<< end >>
