* SPICE3 file created from cmos_inverter.ext - technology: scmos
.include ./ami05.txt
.option scale=0.3u

Vpower vdd gnd 3.3
Vin in gnd PULSE(0 3.3 0 10n 10u 50u 100u)

M1000 out in vdd vdd pfet w=19 l=2
+  ad=95 pd=48 as=95 ps=48
M1001 out in gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
C0 vdd Gnd 3.37fF

.tran 1u 200u
.end
